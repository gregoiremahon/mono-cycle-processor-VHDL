library ieee;
use ieee.std_logic_1164.all;

entity testbench_banc_registres is
end entity testbench_banc_registres;

architecture default of testbench_banc_registres is
    signal clk, rst: std_logic;
    signal w: std_logic_vector(31 downto 0) := (others => '0');
    signal ra, rb, rw: std_logic_vector(3 downto 0) := (others => '0');
    signal we: std_logic := '0';
    signal a, b: std_logic_vector(31 downto 0);

begin
    T0 : entity work.banc_registres
         port map (
             clk => clk,
             rst => rst,
             w => w,
             ra => ra,
             rb => rb,
             rw => rw,
             we => we,
             a => a,
             b => b
         );

    clk_gen : process
    begin
        clk <= '1';
        wait for 2 ns;
        clk <= '0';
        wait for 2 ns;
    end process;

    test : process
    begin
        -- Initialize bank with a reset
        rst <= '1';
        wait for 4 ns;
        rst <= '0';

        -- Read registers @RA = 0 & @RB = 12
        ra <= X"0";
        rb <= X"C";
        -- Wait till values are stabilized
        wait for 1 ns;
        -- Check that we read 0 on both registers
        assert a = X"00000000" report "Error: a is wrong during first read" severity error;
        assert b = X"00000000" report "Error: b is wrong during first read" severity error;

        -- Write into registers @RW = 0 & @RW = 12
        w <= X"0000000A";
        rw <= X"0";
        we <= '1';
        -- Wait for rising edge to pass
        wait for 4 ns;
        rw <= X"C";
        -- Wait for rising edge to pass
        wait for 4 ns;
        we <= '0';

        -- Check that we have successfully written on registers
        ra <= X"0";
        rb <= X"C";
        -- Wait till values are stabilized
        wait for 1 ns;
        -- Check that we read 0xA on both registers
        assert a = X"0000000A" report "Error: a is wrong during second read" severity error;
        assert b = X"0000000A" report "Error: b is wrong during second read" severity error;

        wait;
    end process;

end architecture;

