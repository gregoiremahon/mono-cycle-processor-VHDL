library ieee;
use ieee.std_logic_1164.all;

entity testbench_processing_unit is
end testbench_processing_unit;

architecture arcTB_Processing_Unit of testbench_processing_unit is

    -- Component declaration for the Unit Under Test (UUT)
    component processingUnit
    port (
        clk, rst: in std_logic;
        instruction: in std_logic_vector(31 downto 0);
        dataOut: out std_logic_vector(31 downto 0)
    );
    end component;

    --Inputs
    signal clk : std_logic := '0';
    signal rst : std_logic := '0';
    signal instruction : std_logic_vector(31 downto 0) := (others => '0');

    --Outputs
    signal dataOut : std_logic_vector(31 downto 0);

    -- Clock period definitions
    constant clk_period : time := 10 ns;

begin

    -- Instantiate the Unit Under Test (UUT)
    uut: processingUnit port map (
        clk => clk,
        rst => rst,
        instruction => instruction,
        dataOut => dataOut
    );

    -- Clock process definitions
    clk_process :process
    begin
        clk <= '0';
        wait for clk_period/2;
        clk <= '1';
        wait for clk_period/2;
    end process;

    -- Stimulus process
    stim_proc: process
    begin
        wait for clk_period;

        -- Testcase 1: R(1) = R(15)
        instruction <= "00100000000111110000000000000000"; -- li $15, 42
        wait for clk_period;
        instruction <= "00000000000011110000000100000000"; -- addi $1, $15, 0
        wait for clk_period;
        assert dataOut = x"0000002A" -- 42
        report "Testcase 1 failed" severity error;

        -- Testcase 2: R(1) = R(1) + R(15)
        instruction <= "00100000000111110000000000000000"; -- li $15, 42
        wait for clk_period;
        instruction <= "00000011111000010000000100000000"; -- add $1, $1, $15
        wait for clk_period;
        assert dataOut = x"00000054" -- 42 + 42 = 84
        report "Testcase 2 failed" severity error;
-- Testcase 3: R(2) = R(1) + R(15)
    instruction <= "00100000000111110000000000000000"; -- li $15, 42
    wait for clk_period;
    instruction <= "00000011111000100000001000000000"; -- add $2, $1, $15
    wait for clk_period;
    assert dataOut = x"00000054" -- 42 + 42 = 84
    report "Testcase 3 failed" severity error;

    -- Testcase 4: R(3) = R(1) ? R(15)
    instruction <= "00100000000111110000000000000000"; -- li $15, 42
    wait for clk_period;
    instruction <= "00000011111000110000001100000000"; -- sub $3, $1, $15
    wait for clk_period;
    assert dataOut = x"FFFFFFD6" -- 0 - 42 = -42 (2's complement)
    report "Testcase 4 failed" severity error;

    -- Testcase 5: R(5) = R(7) ? R(15)
    instruction <= "00100000000111110000000000000000"; -- li $15, 42
    wait for clk_period;
    instruction <= "00000111110001100000101100000000"; -- sub $5, $7, $15
    wait for clk_period;
    assert dataOut = x"FFFFFFD6" -- 0 - 42 = -42 (2's complement)
    report "Testcase 5 failed" severity error;

    wait;
end process stim_proc;
end architecture;
